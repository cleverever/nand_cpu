`define PC_SIZE 16
`define BTB_PC_BITS 8
`define CACHE_BLOCK_SIZE 256
`define MEM_TRANS_SIZE 64

import nand_cpu_pkg::*;