module mem_pipeline
(
    
);

endmodule