`define PC_SIZE 16