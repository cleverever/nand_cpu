`define NUM_D_REG 32
`define NUM_S_REG 8

`define PC_SIZE 16
`define BTB_PC_BITS 8
`define CACHE_BLOCK_SIZE 256
`define MEM_TRANS_SIZE 64

`define EX_B_LENGTH 16
`define BR_B_LENGTH 4
`define ST_B_LENGTH 8
`define LD_B_LENGTH 8

`define ROB_LENGTH 64

import nand_cpu_pkg::*;