module nand_cpu
(
    input logic clk,
    input logic n_rst,

    output logic halt
);


//====================================================================================================
//FETCH
//====================================================================================================
fetch_unit FETCH_UNIT();
branch_predictor BRANCH_PREDICTOR();

//----------------------------------------------------------------------------------------------------
//F2D
//----------------------------------------------------------------------------------------------------
fetch_glue FETCH_GLUE();
pr_f2d PR_F2D();

//====================================================================================================
//DECODE
//====================================================================================================
decoder DECODER();
free_list FREE_LIST();
reg_alloc_table REG_ALLOC_TABLE();

//----------------------------------------------------------------------------------------------------
//D2I
//----------------------------------------------------------------------------------------------------
decode_glue DECODE_GLUE();

//====================================================================================================
//ISSUE
//====================================================================================================
regfile REGFILE();

//----------------------------------------------------------------------------------------------------
//I2A
//----------------------------------------------------------------------------------------------------

//====================================================================================================
//ACTION
//====================================================================================================
alu ALU();
d_cache D_CACHE();

//----------------------------------------------------------------------------------------------------
//A2C
//----------------------------------------------------------------------------------------------------

//====================================================================================================
//COMMIT
//====================================================================================================
active_list ACTIVE_LIST();

//XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX
//HAZARD
//XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX
hazard_unit HAZARD_UNIT();

//MMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMMM
//MEMORY
//WWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWWW
memory MEMORY();

endmodule