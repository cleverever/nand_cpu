`include "nand_cpu.svh"

module nand_cpu
(
    input logic clk,
    input logic n_rst,

    output logic halt
);

logic reg_write;
logic [$clog2(`NUM_REG)-1:0] w_addr;

logic p_reg;

logic reg_commit;
logic [$clog2(`NUM_REG)-1:0] commit_addr;

translation_table_ifc translation_table();


//EXECUTION
regfile_ex_ifc ex_rf_read();

//MEMORY

//BRANCH

fetch_unit FETCH_UNIT
(
    .clk,
    .n_rst,

    .interrupt_handler(),

    .i_fetch_ctrl(fetch_ctrl),

    .pc(pc),
    .halted(halt)
);

i_cache I_CACHE
(
    .clk,
    .n_rst,

    .pc(pc),

    .out(f_i_cache_output),

    .cache_request(f_i_cache_request)
);

branch_predictor BRANCH_PREDICTOR
(
    .clk,
    .n_rst,
    
    .pc(pc),

    .use_ps(predictor_use_ps),
    .ps(d_regfile_output.ps),
    
    .out(f_branch_prediction),

    .feedback_valid(a_pr_pass.valid & (a_branch_feedback.branch | a_branch_feedback.jump)),
    .i_feedback(a_branch_feedback)
);

decoder DECODER
(
    .instr(d_instr),
    
    .out(d_decoder_output)
);

free_reg_list FRL
(
    .clk,
    .n_rst,

    .checkin(reg_commit),
    .in(commit_addr),

    .checkout(reg_write),
    .out(p_reg)
);

logic [$clog2(`NUM_REG)-1 : 0] translation [16];

translation_table TT
(
    .clk,
    .n_rst,

    .d_set(reg_write),
    .d_v_reg(w_addr),
    .d_p_reg(p_reg),
    .d_translation(translation)

    .s_set(),
    .s_v_reg(),
    .s_p_reg(),
    .s_translation()
);

regfile RF
(
    .ex_read_request(ex_rf_read),

    .ex_d_write_request(ex_d_write),
    .ex_s_write_request(ex_s_write)
);

execution_buffer EB
(
    .out(execution_buffer_port)
);

e_read_glue E_READ_GLUE
(
    .eb_in(execution_buffer_port),

    .rf_port(ex_rf_read),

    .metadata(e_r_metadata),
    .rf_dst(e_r_rf_dst),
    .alu_input(r_alu_input)
);

metadata_ifc e_r_metadata();
rf_dst_ifc e_r_rf_dst();
alu_input_ifc r_alu_input();

e_r2a E_R2A
(
    .md_in(e_r_metadata),
    .rf_dst_in(e_r_rf_dst),
    .alu_input_in(r_alu_input),

    .md_out(e_a_metadata),
    .rf_dst_out(e_a_rf_dst),
    .alu_input_out(a_alu_input)
);

metadata_ifc e_a_metadata();
rf_dst_ifc e_a_rf_dst();
alu_input_ifc a_alu_input();

alu ALU
(
    .in(a_alu_input),
    .out(alu_output)
);

logic [15:0] alu_output;

e_alu_glue E_ALU_GLUE
(
    .alu_result(alu_output),

    .ex_d_write(e_a_d_write),
    .ex_s_write(e_a_s_write)
);

regfile_d_write_ifc e_a_d_write();
regfile_s_write_ifc e_a_s_write();

e_a2c E_A2C
(
    .md_in(e_a_metadata),
    .e_a_d_write(e_a_d_write),
    .e_a_s_write(e_a_s_write),

    .md_out(e_c_metadata),
    .e_c_d_write(ex_d_write),
    .e_c_s_write(ex_s_write)
);

metadata_ifc e_c_metadata();
regfile_d_write_ifc ex_d_write();
regfile_s_write_ifc ex_s_write();

reorder_buffer ROB
(
    .reg_write(reg_commit),
    .reg_addr(commit_addr)
);

endmodule