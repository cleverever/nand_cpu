module ar_pipeline
(
    
);

endmodule