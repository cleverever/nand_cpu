`define PC_SIZE 16

import nand_cpu_pkg::*;