`define DATA_WIDTH 16
`define NUM_REG 16