`define PC_SIZE 16
`define BTB_PC_BITS 8

import nand_cpu_pkg::*;