`define PC_SIZE 16
`define NUM_REG 32
`define NUM_PS 2
`define AL_SIZE 20

import nand_cpu_pkg::*;